	sbox0[0] = 14;
	sbox0[1] = 0;
	sbox0[2] = 4;
	sbox0[3] = 15;
	sbox0[4] = 13;
	sbox0[5] = 7;
	sbox0[6] = 1;
	sbox0[7] = 4;
	sbox0[8] = 2;
	sbox0[9] = 14;
	sbox0[10] = 15;
	sbox0[11] = 2;
	sbox0[12] = 11;
	sbox0[13] = 13;
	sbox0[14] = 8;
	sbox0[15] = 1;
	sbox0[16] = 3;
	sbox0[17] = 10;
	sbox0[18] = 10;
	sbox0[19] = 6;
	sbox0[20] = 6;
	sbox0[21] = 12;
	sbox0[22] = 12;
	sbox0[23] = 11;
	sbox0[24] = 5;
	sbox0[25] = 9;
	sbox0[26] = 9;
	sbox0[27] = 5;
	sbox0[28] = 0;
	sbox0[29] = 3;
	sbox0[30] = 7;
	sbox0[31] = 8;
	sbox0[32] = 4;
	sbox0[33] = 15;
	sbox0[34] = 1;
	sbox0[35] = 12;
	sbox0[36] = 14;
	sbox0[37] = 8;
	sbox0[38] = 8;
	sbox0[39] = 2;
	sbox0[40] = 13;
	sbox0[41] = 4;
	sbox0[42] = 6;
	sbox0[43] = 9;
	sbox0[44] = 2;
	sbox0[45] = 1;
	sbox0[46] = 11;
	sbox0[47] = 7;
	sbox0[48] = 15;
	sbox0[49] = 5;
	sbox0[50] = 12;
	sbox0[51] = 11;
	sbox0[52] = 9;
	sbox0[53] = 3;
	sbox0[54] = 7;
	sbox0[55] = 14;
	sbox0[56] = 3;
	sbox0[57] = 10;
	sbox0[58] = 10;
	sbox0[59] = 0;
	sbox0[60] = 5;
	sbox0[61] = 6;
	sbox0[62] = 0;
	sbox0[63] = 13;
	sbox1[0] = 15;
	sbox1[1] = 3;
	sbox1[2] = 1;
	sbox1[3] = 13;
	sbox1[4] = 8;
	sbox1[5] = 4;
	sbox1[6] = 14;
	sbox1[7] = 7;
	sbox1[8] = 6;
	sbox1[9] = 15;
	sbox1[10] = 11;
	sbox1[11] = 2;
	sbox1[12] = 3;
	sbox1[13] = 8;
	sbox1[14] = 4;
	sbox1[15] = 14;
	sbox1[16] = 9;
	sbox1[17] = 12;
	sbox1[18] = 7;
	sbox1[19] = 0;
	sbox1[20] = 2;
	sbox1[21] = 1;
	sbox1[22] = 13;
	sbox1[23] = 10;
	sbox1[24] = 12;
	sbox1[25] = 6;
	sbox1[26] = 0;
	sbox1[27] = 9;
	sbox1[28] = 5;
	sbox1[29] = 11;
	sbox1[30] = 10;
	sbox1[31] = 5;
	sbox1[32] = 0;
	sbox1[33] = 13;
	sbox1[34] = 14;
	sbox1[35] = 8;
	sbox1[36] = 7;
	sbox1[37] = 10;
	sbox1[38] = 11;
	sbox1[39] = 1;
	sbox1[40] = 10;
	sbox1[41] = 3;
	sbox1[42] = 4;
	sbox1[43] = 15;
	sbox1[44] = 13;
	sbox1[45] = 4;
	sbox1[46] = 1;
	sbox1[47] = 2;
	sbox1[48] = 5;
	sbox1[49] = 11;
	sbox1[50] = 8;
	sbox1[51] = 6;
	sbox1[52] = 12;
	sbox1[53] = 7;
	sbox1[54] = 6;
	sbox1[55] = 12;
	sbox1[56] = 9;
	sbox1[57] = 0;
	sbox1[58] = 3;
	sbox1[59] = 5;
	sbox1[60] = 2;
	sbox1[61] = 14;
	sbox1[62] = 15;
	sbox1[63] = 9;
	sbox2[0] = 10;
	sbox2[1] = 13;
	sbox2[2] = 0;
	sbox2[3] = 7;
	sbox2[4] = 9;
	sbox2[5] = 0;
	sbox2[6] = 14;
	sbox2[7] = 9;
	sbox2[8] = 6;
	sbox2[9] = 3;
	sbox2[10] = 3;
	sbox2[11] = 4;
	sbox2[12] = 15;
	sbox2[13] = 6;
	sbox2[14] = 5;
	sbox2[15] = 10;
	sbox2[16] = 1;
	sbox2[17] = 2;
	sbox2[18] = 13;
	sbox2[19] = 8;
	sbox2[20] = 12;
	sbox2[21] = 5;
	sbox2[22] = 7;
	sbox2[23] = 14;
	sbox2[24] = 11;
	sbox2[25] = 12;
	sbox2[26] = 4;
	sbox2[27] = 11;
	sbox2[28] = 2;
	sbox2[29] = 15;
	sbox2[30] = 8;
	sbox2[31] = 1;
	sbox2[32] = 13;
	sbox2[33] = 1;
	sbox2[34] = 6;
	sbox2[35] = 10;
	sbox2[36] = 4;
	sbox2[37] = 13;
	sbox2[38] = 9;
	sbox2[39] = 0;
	sbox2[40] = 8;
	sbox2[41] = 6;
	sbox2[42] = 15;
	sbox2[43] = 9;
	sbox2[44] = 3;
	sbox2[45] = 8;
	sbox2[46] = 0;
	sbox2[47] = 7;
	sbox2[48] = 11;
	sbox2[49] = 4;
	sbox2[50] = 1;
	sbox2[51] = 15;
	sbox2[52] = 2;
	sbox2[53] = 14;
	sbox2[54] = 12;
	sbox2[55] = 3;
	sbox2[56] = 5;
	sbox2[57] = 11;
	sbox2[58] = 10;
	sbox2[59] = 5;
	sbox2[60] = 14;
	sbox2[61] = 2;
	sbox2[62] = 7;
	sbox2[63] = 12;
	sbox3[0] = 7;
	sbox3[1] = 13;
	sbox3[2] = 13;
	sbox3[3] = 8;
	sbox3[4] = 14;
	sbox3[5] = 11;
	sbox3[6] = 3;
	sbox3[7] = 5;
	sbox3[8] = 0;
	sbox3[9] = 6;
	sbox3[10] = 6;
	sbox3[11] = 15;
	sbox3[12] = 9;
	sbox3[13] = 0;
	sbox3[14] = 10;
	sbox3[15] = 3;
	sbox3[16] = 1;
	sbox3[17] = 4;
	sbox3[18] = 2;
	sbox3[19] = 7;
	sbox3[20] = 8;
	sbox3[21] = 2;
	sbox3[22] = 5;
	sbox3[23] = 12;
	sbox3[24] = 11;
	sbox3[25] = 1;
	sbox3[26] = 12;
	sbox3[27] = 10;
	sbox3[28] = 4;
	sbox3[29] = 14;
	sbox3[30] = 15;
	sbox3[31] = 9;
	sbox3[32] = 10;
	sbox3[33] = 3;
	sbox3[34] = 6;
	sbox3[35] = 15;
	sbox3[36] = 9;
	sbox3[37] = 0;
	sbox3[38] = 0;
	sbox3[39] = 6;
	sbox3[40] = 12;
	sbox3[41] = 10;
	sbox3[42] = 11;
	sbox3[43] = 1;
	sbox3[44] = 7;
	sbox3[45] = 13;
	sbox3[46] = 13;
	sbox3[47] = 8;
	sbox3[48] = 15;
	sbox3[49] = 9;
	sbox3[50] = 1;
	sbox3[51] = 4;
	sbox3[52] = 3;
	sbox3[53] = 5;
	sbox3[54] = 14;
	sbox3[55] = 11;
	sbox3[56] = 5;
	sbox3[57] = 12;
	sbox3[58] = 2;
	sbox3[59] = 7;
	sbox3[60] = 8;
	sbox3[61] = 2;
	sbox3[62] = 4;
	sbox3[63] = 14;
	sbox4[0] = 2;
	sbox4[1] = 14;
	sbox4[2] = 12;
	sbox4[3] = 11;
	sbox4[4] = 4;
	sbox4[5] = 2;
	sbox4[6] = 1;
	sbox4[7] = 12;
	sbox4[8] = 7;
	sbox4[9] = 4;
	sbox4[10] = 10;
	sbox4[11] = 7;
	sbox4[12] = 11;
	sbox4[13] = 13;
	sbox4[14] = 6;
	sbox4[15] = 1;
	sbox4[16] = 8;
	sbox4[17] = 5;
	sbox4[18] = 5;
	sbox4[19] = 0;
	sbox4[20] = 3;
	sbox4[21] = 15;
	sbox4[22] = 15;
	sbox4[23] = 10;
	sbox4[24] = 13;
	sbox4[25] = 3;
	sbox4[26] = 0;
	sbox4[27] = 9;
	sbox4[28] = 14;
	sbox4[29] = 8;
	sbox4[30] = 9;
	sbox4[31] = 6;
	sbox4[32] = 4;
	sbox4[33] = 11;
	sbox4[34] = 2;
	sbox4[35] = 8;
	sbox4[36] = 1;
	sbox4[37] = 12;
	sbox4[38] = 11;
	sbox4[39] = 7;
	sbox4[40] = 10;
	sbox4[41] = 1;
	sbox4[42] = 13;
	sbox4[43] = 14;
	sbox4[44] = 7;
	sbox4[45] = 2;
	sbox4[46] = 8;
	sbox4[47] = 13;
	sbox4[48] = 15;
	sbox4[49] = 6;
	sbox4[50] = 9;
	sbox4[51] = 15;
	sbox4[52] = 12;
	sbox4[53] = 0;
	sbox4[54] = 5;
	sbox4[55] = 9;
	sbox4[56] = 6;
	sbox4[57] = 10;
	sbox4[58] = 3;
	sbox4[59] = 4;
	sbox4[60] = 0;
	sbox4[61] = 5;
	sbox4[62] = 14;
	sbox4[63] = 3;
	sbox5[0] = 12;
	sbox5[1] = 10;
	sbox5[2] = 1;
	sbox5[3] = 15;
	sbox5[4] = 10;
	sbox5[5] = 4;
	sbox5[6] = 15;
	sbox5[7] = 2;
	sbox5[8] = 9;
	sbox5[9] = 7;
	sbox5[10] = 2;
	sbox5[11] = 12;
	sbox5[12] = 6;
	sbox5[13] = 9;
	sbox5[14] = 8;
	sbox5[15] = 5;
	sbox5[16] = 0;
	sbox5[17] = 6;
	sbox5[18] = 13;
	sbox5[19] = 1;
	sbox5[20] = 3;
	sbox5[21] = 13;
	sbox5[22] = 4;
	sbox5[23] = 14;
	sbox5[24] = 14;
	sbox5[25] = 0;
	sbox5[26] = 7;
	sbox5[27] = 11;
	sbox5[28] = 5;
	sbox5[29] = 3;
	sbox5[30] = 11;
	sbox5[31] = 8;
	sbox5[32] = 9;
	sbox5[33] = 4;
	sbox5[34] = 14;
	sbox5[35] = 3;
	sbox5[36] = 15;
	sbox5[37] = 2;
	sbox5[38] = 5;
	sbox5[39] = 12;
	sbox5[40] = 2;
	sbox5[41] = 9;
	sbox5[42] = 8;
	sbox5[43] = 5;
	sbox5[44] = 12;
	sbox5[45] = 15;
	sbox5[46] = 3;
	sbox5[47] = 10;
	sbox5[48] = 7;
	sbox5[49] = 11;
	sbox5[50] = 0;
	sbox5[51] = 14;
	sbox5[52] = 4;
	sbox5[53] = 1;
	sbox5[54] = 10;
	sbox5[55] = 7;
	sbox5[56] = 1;
	sbox5[57] = 6;
	sbox5[58] = 13;
	sbox5[59] = 0;
	sbox5[60] = 11;
	sbox5[61] = 8;
	sbox5[62] = 6;
	sbox5[63] = 13;
	sbox6[0] = 4;
	sbox6[1] = 13;
	sbox6[2] = 11;
	sbox6[3] = 0;
	sbox6[4] = 2;
	sbox6[5] = 11;
	sbox6[6] = 14;
	sbox6[7] = 7;
	sbox6[8] = 15;
	sbox6[9] = 4;
	sbox6[10] = 0;
	sbox6[11] = 9;
	sbox6[12] = 8;
	sbox6[13] = 1;
	sbox6[14] = 13;
	sbox6[15] = 10;
	sbox6[16] = 3;
	sbox6[17] = 14;
	sbox6[18] = 12;
	sbox6[19] = 3;
	sbox6[20] = 9;
	sbox6[21] = 5;
	sbox6[22] = 7;
	sbox6[23] = 12;
	sbox6[24] = 5;
	sbox6[25] = 2;
	sbox6[26] = 10;
	sbox6[27] = 15;
	sbox6[28] = 6;
	sbox6[29] = 8;
	sbox6[30] = 1;
	sbox6[31] = 6;
	sbox6[32] = 1;
	sbox6[33] = 6;
	sbox6[34] = 4;
	sbox6[35] = 11;
	sbox6[36] = 11;
	sbox6[37] = 13;
	sbox6[38] = 13;
	sbox6[39] = 8;
	sbox6[40] = 12;
	sbox6[41] = 1;
	sbox6[42] = 3;
	sbox6[43] = 4;
	sbox6[44] = 7;
	sbox6[45] = 10;
	sbox6[46] = 14;
	sbox6[47] = 7;
	sbox6[48] = 10;
	sbox6[49] = 9;
	sbox6[50] = 15;
	sbox6[51] = 5;
	sbox6[52] = 6;
	sbox6[53] = 0;
	sbox6[54] = 8;
	sbox6[55] = 15;
	sbox6[56] = 0;
	sbox6[57] = 14;
	sbox6[58] = 5;
	sbox6[59] = 2;
	sbox6[60] = 9;
	sbox6[61] = 3;
	sbox6[62] = 2;
	sbox6[63] = 12;
	sbox7[0] = 13;
	sbox7[1] = 1;
	sbox7[2] = 2;
	sbox7[3] = 15;
	sbox7[4] = 8;
	sbox7[5] = 13;
	sbox7[6] = 4;
	sbox7[7] = 8;
	sbox7[8] = 6;
	sbox7[9] = 10;
	sbox7[10] = 15;
	sbox7[11] = 3;
	sbox7[12] = 11;
	sbox7[13] = 7;
	sbox7[14] = 1;
	sbox7[15] = 4;
	sbox7[16] = 10;
	sbox7[17] = 12;
	sbox7[18] = 9;
	sbox7[19] = 5;
	sbox7[20] = 3;
	sbox7[21] = 6;
	sbox7[22] = 14;
	sbox7[23] = 11;
	sbox7[24] = 5;
	sbox7[25] = 0;
	sbox7[26] = 0;
	sbox7[27] = 14;
	sbox7[28] = 12;
	sbox7[29] = 9;
	sbox7[30] = 7;
	sbox7[31] = 2;
	sbox7[32] = 7;
	sbox7[33] = 2;
	sbox7[34] = 11;
	sbox7[35] = 1;
	sbox7[36] = 4;
	sbox7[37] = 14;
	sbox7[38] = 1;
	sbox7[39] = 7;
	sbox7[40] = 9;
	sbox7[41] = 4;
	sbox7[42] = 12;
	sbox7[43] = 10;
	sbox7[44] = 14;
	sbox7[45] = 8;
	sbox7[46] = 2;
	sbox7[47] = 13;
	sbox7[48] = 0;
	sbox7[49] = 15;
	sbox7[50] = 6;
	sbox7[51] = 12;
	sbox7[52] = 10;
	sbox7[53] = 9;
	sbox7[54] = 13;
	sbox7[55] = 0;
	sbox7[56] = 15;
	sbox7[57] = 3;
	sbox7[58] = 3;
	sbox7[59] = 5;
	sbox7[60] = 5;
	sbox7[61] = 6;
	sbox7[62] = 8;
	sbox7[63] = 11;
